* /home/drako/eSim-Workspace/xor_gate/xor_gate.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jun 29 19:54:09 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M3  Net-_M13-Pad2_ /b Net-_M3-Pad3_ Net-_M3-Pad3_ mosfet_n		
M6  Net-_M5-Pad3_ Net-_M11-Pad3_ Net-_M13-Pad2_ Net-_M5-Pad3_ mosfet_p		
M5  Net-_M11-Pad1_ /b Net-_M5-Pad3_ Net-_M11-Pad1_ mosfet_p		
M8  Net-_M5-Pad3_ /a Net-_M13-Pad2_ Net-_M5-Pad3_ mosfet_p		
M4  Net-_M3-Pad3_ Net-_M1-Pad1_ GND GND mosfet_n		
M9  Net-_M13-Pad2_ Net-_M11-Pad3_ Net-_M10-Pad1_ Net-_M10-Pad1_ mosfet_n		
M10  Net-_M10-Pad1_ /a GND GND mosfet_n		
M12  Net-_M11-Pad3_ /b GND GND mosfet_n		
M11  Net-_M11-Pad1_ /b Net-_M11-Pad3_ Net-_M11-Pad1_ mosfet_p		
M1  Net-_M1-Pad1_ /a GND GND mosfet_n		
M2  Net-_M11-Pad1_ /a Net-_M1-Pad1_ Net-_M11-Pad1_ mosfet_p		
U1  /a /b /yout PORT		
M13  /yout Net-_M13-Pad2_ GND GND mosfet_n		
M14  Net-_M11-Pad1_ Net-_M13-Pad2_ /yout Net-_M11-Pad1_ mosfet_p		
M7  Net-_M11-Pad1_ Net-_M1-Pad1_ Net-_M5-Pad3_ Net-_M11-Pad1_ mosfet_p		
v1  Net-_M11-Pad1_ GND 3.3v		

.end
