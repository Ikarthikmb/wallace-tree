* /home/drako/eSim-Workspace/halfadder/halfadder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jun 29 20:24:42 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  /CARRY /SUM PORT		
U2  /a0 /b0 PORT		
x2  /a0 /b0 /CARRY and_gate		
x1  /a0 /b0 /SUM xor_gate		

.end
