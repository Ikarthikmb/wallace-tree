* /home/drako/applications/esim-2.1/library/subcircuitlibrary/and_gate/and_gate.cir

.lib "~/eSim-Workspace/prelayout/sky130_fd_pr/models/sky130.lib.spice" tt

xm2  net-_m1-pad3_ a net-_m2-pad3_ net-_m2-pad3_ sky130_fd_pr__nfet_01v8 w=1 l=0.5 m=1
xm3  net-_m2-pad3_ b gnd gnd sky130_fd_pr__nfet_01v8 w=1 l=0.5 m=1
xm1  vdd a net-_m1-pad3_ vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5 m=1
xm4  vdd b net-_m1-pad3_ vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5 m=1
xm5  out net-_m1-pad3_ gnd gnd sky130_fd_pr__nfet_01v8 w=1 l=0.5 m=1
xm6  vdd net-_m1-pad3_ out vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5 m=1
* u1  a b out port
v1 vdd gnd  dc 3.3
.tran 0e-00 0e-00 0e-00

* Control Statements 
.control
run
print allv > plot_data_v.txt
print alli > plot_data_i.txt
.endc
.end
