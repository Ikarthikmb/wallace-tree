* /home/drako/esim-workspace/wallace3tree/wallace3tree.cir

.lib "~/eSim-Workspace/prelayout/sky130_fd_pr/models/sky130.lib.spice" tt

.include fulladder.sub
.include and_gate.sub
.include halfadder.sub
x2 b0 a0 z0 and_gate
x1 b0 a1 net-_x1-pad3_ and_gate
x5 b1 a0 net-_x5-pad3_ and_gate
x6 b1 a1 net-_x6-pad3_ and_gate
x7 net-_x5-pad3_ net-_x1-pad3_ z1 net-_x7-pad4_ halfadder
* u1  a1 a0 a2 b0 b1 b2 z0 z1 z2 z3 z4 z5 port
x3 b0 a2 net-_x3-pad3_ and_gate
x4 b1 a2 net-_x4-pad3_ and_gate
x8 net-_x6-pad3_ net-_x3-pad3_ net-_x7-pad4_ net-_x13-pad2_ net-_x8-pad5_ fulladder
x10 b2 a0 net-_x10-pad3_ and_gate
x11 b2 a1 net-_x11-pad3_ and_gate
x12 b2 a2 net-_x12-pad3_ and_gate
x13 net-_x10-pad3_ net-_x13-pad2_ z2 net-_x13-pad4_ halfadder
x14 net-_x11-pad3_ net-_x14-pad2_ net-_x13-pad4_ z3 net-_x14-pad5_ fulladder
x9 net-_x8-pad5_ net-_x4-pad3_ net-_x14-pad2_ net-_x15-pad2_ halfadder
x15 net-_x12-pad3_ net-_x15-pad2_ net-_x14-pad5_ z4 z5 fulladder

v1 a0 0 pulse 0 1.8 0 0 0 5m 10m
v2 a1 0 pulse 0 1.8 10m 0 0 5m 15m
v3 a2 0 pulse 0 1.8 0 0 0 5m 10m

v4 b0 0 pulse 0 1.8 5m 0 0 5m 10m
v5 b1 0 pulse 0 1.8 0 0 0 15m 30m
v6 b2 0 pulse 0 1.8 10m 0 0 5m 15m

.tran 0.1m 20m

* Control Statements 
.control
run
plot a0
plot a1
plot a2
plot b0
plot b1
plot b2

plot z0
plot z1
plot z2
plot z3
plot z4
plot z5

print allv > plot_data_v.txt
print alli > plot_data_i.txt
.endc
.end
